interface clock_if;

    logic clock;

endinterface: clock_if
