package test_clock;
    
    import uvm_pkg::*;

    `include "env_config.svh"
    `include "env.svh"
    `include "test.svh"


endpackage: test_clock